--------------------------------------------------------------------------------
-- Title         : 3-bit Comparator
-- Project       : VHDL Synthesis Overview
-------------------------------------------------------------------------------
-- File          : threeBitComparator.vhd
-- Author        : Rami Abielmona  <rabielmo@site.uottawa.ca>
-- Created       : 2003/05/17
-- Last modified : 2007/09/25
-------------------------------------------------------------------------------
-- Description : This file creates a 3-bit binary comparator as defined in the VHDL
--		 Synthesis lecture.  The architecture is done at the RTL
--		 abstraction level and the implementation is done in structural
--		 VHDL.
-------------------------------------------------------------------------------
-- Modification history :
-- 2003.05.17 	R. Abielmona		Creation
-- 2004.09.22 	R. Abielmona		Ported for CEG 3550
-- 2007.09.25 	R. Abielmona		Modified copyright notice
-------------------------------------------------------------------------------
-- This file is copyright material of Rami Abielmona, Ph.D., P.Eng., Chief Research
-- Scientist at Larus Technologies.  Permission to make digital or hard copies of part
-- or all of this work for personal or classroom use is granted without fee
-- provided that copies are not made or distributed for profit or commercial
-- advantage and that copies bear this notice and the full citation of this work.
-- Prior permission is required to copy, republish, redistribute or post this work.
-- This notice is adapted from the ACM copyright notice.
--------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY fourBitComparator IS
    PORT(
        i_Ai, i_Bi : IN  STD_LOGIC_VECTOR(3 downto 0);
        o_GT, o_LT, o_EQ : OUT STD_LOGIC
    );
END fourBitComparator;

ARCHITECTURE rtl OF fourBitComparator IS
    SIGNAL int_GT, int_LT : STD_LOGIC_VECTOR(3 downto 0);
    SIGNAL gnd : STD_LOGIC;

    COMPONENT oneBitComparator
        PORT(
            i_GTPrevious, i_LTPrevious : IN  STD_LOGIC;
            i_Ai, i_Bi : IN  STD_LOGIC;
            o_GT, o_LT : OUT STD_LOGIC
        );
    END COMPONENT;
BEGIN
    -- Concurrent Signal Assignment
    gnd <= '0';

    comp3: oneBitComparator
        PORT MAP (
            i_GTPrevious => gnd,
            i_LTPrevious => gnd,
            i_Ai => i_Ai(3),
            i_Bi => i_Bi(3),
            o_GT => int_GT(3),
            o_LT => int_LT(3)
        );

    comp2: oneBitComparator
        PORT MAP (
            i_GTPrevious => int_GT(3),
            i_LTPrevious => int_LT(3),
            i_Ai => i_Ai(2),
            i_Bi => i_Bi(2),
            o_GT => int_GT(2),
            o_LT => int_LT(2)
        );

    comp1: oneBitComparator
        PORT MAP (
            i_GTPrevious => int_GT(2),
            i_LTPrevious => int_LT(2),
            i_Ai => i_Ai(1),
            i_Bi => i_Bi(1),
            o_GT => int_GT(1),
            o_LT => int_LT(1)
        );

    comp0: oneBitComparator
        PORT MAP (
            i_GTPrevious => int_GT(1),
            i_LTPrevious => int_LT(1),
            i_Ai => i_Ai(0),
            i_Bi => i_Bi(0),
            o_GT => int_GT(0),
            o_LT => int_LT(0)
        );

    -- Output Driver
    o_GT <= int_GT(0);
    o_LT <= int_LT(0);
    o_EQ <= int_GT(0) nor int_LT(0);

END rtl;
