LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY fourBitRegister_Counter IS
  PORT (
    i_resetBar : IN  STD_LOGIC;                       -- async reset, active low
    i_clock    : IN  STD_LOGIC;
    i_sel_0    : IN  STD_LOGIC;                       -- control select (LSB)
    i_sel_1    : IN  STD_LOGIC;                       -- control select (MSB)
    i_Value    : IN  STD_LOGIC_VECTOR(3 downto 0);    -- parallel load value
    o_Value    : OUT STD_LOGIC_VECTOR(3 downto 0);    -- register contents
    o_zero     : OUT STD_LOGIC                        -- flag when value=0000
  );
END fourBitRegister_Counter;

ARCHITECTURE rtl OF fourBitRegister_Counter IS
  SIGNAL int_Value : STD_LOGIC_VECTOR(3 downto 0);  -- Q (current)
  SIGNAL inc_Value : STD_LOGIC_VECTOR(3 downto 0);  -- Q + 1
  SIGNAL nxt_Value : STD_LOGIC_VECTOR(3 downto 0);  -- D (next)

  COMPONENT enARdFF_2
    PORT(
      i_resetBar : IN  STD_LOGIC;
      i_d        : IN  STD_LOGIC;
      i_enable   : IN  STD_LOGIC;
      i_clock    : IN  STD_LOGIC;
      o_q        : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT Mux4_1 IS
    PORT(
      i_val_0, i_val_1, i_val_2, i_val_3 : IN STD_LOGIC;
      i_sel_0, i_sel_1 : IN STD_LOGIC;
      o_val : OUT STD_LOGIC
    );
  END COMPONENT;

  -- carry chain for incrementer
  SIGNAL c1, c2, c3 : STD_LOGIC;
BEGIN
  -------------------------------------------------------------------
  -- Ripple-carry incrementer: inc_Value = int_Value + 1 (mod 16)
  -------------------------------------------------------------------
  inc_Value(0) <= NOT int_Value(0);
  c1           <= int_Value(0);

  inc_Value(1) <= int_Value(1) XOR c1;
  c2           <= int_Value(1) AND c1;

  inc_Value(2) <= int_Value(2) XOR c2;
  c3           <= int_Value(2) AND c2;

  inc_Value(3) <= int_Value(3) XOR c3;

  -------------------------------------------------------------------
  -- MUX + FF for each bit
  -- 00: Hold (Q), 01: Load (i_Value), 10: Up, 11: Up
  -------------------------------------------------------------------
  bit3MUX : Mux4_1 PORT MAP(
    i_val_0 => int_Value(3),   -- Hold
    i_val_1 => i_Value(3),     -- Load
    i_val_2 => inc_Value(3),   -- Up
    i_val_3 => inc_Value(3),   -- Up
    i_sel_0 => i_sel_0, i_sel_1 => i_sel_1,
    o_val   => nxt_Value(3)
  );
  bit3FF : enARdFF_2 PORT MAP(i_resetBar=>i_resetBar, i_d=>nxt_Value(3), i_enable=>'1', i_clock=>i_clock, o_q=>int_Value(3));

  bit2MUX : Mux4_1 PORT MAP(
    i_val_0 => int_Value(2),
    i_val_1 => i_Value(2),
    i_val_2 => inc_Value(2),
    i_val_3 => inc_Value(2),
    i_sel_0 => i_sel_0, i_sel_1 => i_sel_1,
    o_val   => nxt_Value(2)
  );
  bit2FF : enARdFF_2 PORT MAP(i_resetBar=>i_resetBar, i_d=>nxt_Value(2), i_enable=>'1', i_clock=>i_clock, o_q=>int_Value(2));

  bit1MUX : Mux4_1 PORT MAP(
    i_val_0 => int_Value(1),
    i_val_1 => i_Value(1),
    i_val_2 => inc_Value(1),
    i_val_3 => inc_Value(1),
    i_sel_0 => i_sel_0, i_sel_1 => i_sel_1,
    o_val   => nxt_Value(1)
  );
  bit1FF : enARdFF_2 PORT MAP(i_resetBar=>i_resetBar, i_d=>nxt_Value(1), i_enable=>'1', i_clock=>i_clock, o_q=>int_Value(1));

  bit0MUX : Mux4_1 PORT MAP(
    i_val_0 => int_Value(0),
    i_val_1 => i_Value(0),
    i_val_2 => inc_Value(0),
    i_val_3 => inc_Value(0),
    i_sel_0 => i_sel_0, i_sel_1 => i_sel_1,
    o_val   => nxt_Value(0)
  );
  bit0FF : enARdFF_2 PORT MAP(i_resetBar=>i_resetBar, i_d=>nxt_Value(0), i_enable=>'1', i_clock=>i_clock, o_q=>int_Value(0));

  -------------------------------------------------------------------
  -- Outputs
  -------------------------------------------------------------------
  o_Value <= int_Value;
  o_zero  <= '1' WHEN int_Value="0000" ELSE '0';
END rtl;
